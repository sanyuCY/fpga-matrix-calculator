`timescale 1ns / 1ps




module control_fsm(
    input clk,                  // ȫ��ʱ�ӣ�100MHz��
    input rst_n,                // ȫ�ָ�λ���͵�ƽ��Ч��
    input [7:0] SW,             // 8λ���뿪�أ�SW0~SW7��
    input [4:0] KEY,            // 5λ������S1~S5��ӦKEY[0]~KEY[4]��
    input op_done,              // ������ɱ�־�����Գ�ԱC��
    input input_done,           // ����/������ɱ�־�����Գ�ԱC��
    input display_done,         // չʾ��ɱ�־�����Գ�ԱA��
    input [2:0] error_type,     // �������ͣ����Գ�ԱC��000=�޴�
    input [7:0] uart_rx_data,   // ����ָ����Գ�ԱA��
    input rx_done,              // ����ָ�������ɣ����Գ�ԱA��
    input [3:0] max_mat_num,    // �������洢����������param_config��
    input [7:0] val_min,        // Ԫ����Сֵ������param_config��
    input [7:0] val_max,        // Ԫ�����ֵ������param_config��
    input config_done,          // ������ɱ�־������param_config��
    input [3:0] result_m,       // ����������������Գ�ԱC��
    input [3:0] result_n,       // ����������������Գ�ԱC��
    output reg [3:0] current_mode,  // ��ǰ״̬�����������ģ�飩
    output reg [2:0] current_op,    // �������ͣ��������ԱC��
    output reg [7:0] LED,           // LED���ƣ�����������壩
    output reg [15:0] seg_code,     // ����ܿ��ƣ�16λ����4+��4��
    output reg [3:0] scalar,        // ����ֵ���������ԱC��
    output reg [1:0] operand_sel,   // ������ѡ��ģʽ��00=�ֶ���01=�����
    output reg [3:0] countdown_sec  // ����ʱ�������������ԱA��
);

// 1. ״̬���壨9������״̬��
localparam S_MENU      = 4'b0000;  // ���˵�
localparam S_INPUT     = 4'b0001;  // ��������ģʽ
localparam S_GEN       = 4'b0010;  // ��������ģʽ
localparam S_SHOW      = 4'b0011;  // ����չʾģʽ
localparam S_OP_SELECT = 4'b0100;  // ѡ����������
localparam S_OP_PARAM  = 4'b0101;  // ѡ��������
localparam S_OP_EXEC   = 4'b0110;  // ִ������
localparam S_RESULT    = 4'b0111;  // չʾ���
localparam S_RETURN    = 4'b1000;  // �ȴ�����

// 2. �������ͱ��루��SW0~SW2��Ӧ��
localparam OP_TRANS    = 3'b000;  // ת�� T
localparam OP_ADD      = 3'b001;  // �ӷ� A
localparam OP_SCALAR   = 3'b010;  // ������ B
localparam OP_MUL      = 3'b011;  // ����� C
localparam OP_CONV     = 3'b100;  // ��� J��bonus��

// 3. �������ʾ���루��������XC7A35T���ݣ�
localparam SEG_OFF     = 8'b11111111;  // Ϩ��
localparam SEG_0       = 8'b00000011;  // 0
localparam SEG_1       = 8'b10011111;  // 1
localparam SEG_2       = 8'b01001001;  // 2
localparam SEG_3       = 8'b01001101;  // 3
localparam SEG_4       = 8'b00100111;  // 4
localparam SEG_5       = 8'b00101101;  // 5
localparam SEG_6       = 8'b00111101;  // 6
localparam SEG_7       = 8'b01000011;  // 7
localparam SEG_8       = 8'b00000001;  // 8
localparam SEG_9       = 8'b00000101;  // 9
localparam SEG_T       = 8'b01010001;  // T
localparam SEG_A       = 8'b00010001;  // A
localparam SEG_B       = 8'b00110001;  // B
localparam SEG_C       = 8'b01000101;  // C
localparam SEG_J       = 8'b01011001;  // J

// 4. ���������ض��壨100MHzʱ�����䣩
reg [23:0] key_cnt;           // ����������������100MHz*10ms=1,000,000��
reg [4:0] key_sync;           // ����ͬ���Ĵ���
reg [4:0] key_clean;          // ������İ����źţ��ߵ�ƽ��Ч��
reg [23:0] sw_cnt;            // ���뿪�ط���������
reg [7:0] sw_sync;            // ���뿪��ͬ���Ĵ���
reg [7:0] sw_clean;           // ������Ĳ��뿪���ź�
reg [31:0] countdown_cnt;     // ���󵹼�ʱ��������100MHzʱ�ӣ�
reg countdown_en;             // ����ʱʹ���ź�
reg [3:0] countdown_cfg;      // ����ʱ����ֵ��5~15�룬Ĭ��10�룩

// 5. ��λ��ʼ�����͵�ƽ��Ч��
always @(negedge rst_n) begin
    current_mode <= S_MENU;       // ��λ��ص����˵�
    current_op <= OP_TRANS;       // Ĭ���������ͣ�ת��
    LED <= 8'b00000000;           // ����LEDϨ��
    seg_code <= {SEG_OFF, SEG_OFF};// �����Ϩ��
    scalar <= 4'd0;               // ����Ĭ��0
    operand_sel <= 2'b00;         // Ĭ���ֶ�ѡ��������
    key_cnt <= 24'd0;
    key_sync <= 5'b00000;
    key_clean <= 5'b00000;
    sw_cnt <= 24'd0;
    sw_sync <= 8'b00000000;
    sw_clean <= 8'b00000000;
    countdown_cnt <= 32'd0;
    countdown_sec <= 4'd10;       // Ĭ�ϵ���ʱ10��
    countdown_cfg <= 4'd10;       // Ĭ������10��
    countdown_en <= 1'b0;
end

// 6. ���������߼���100MHzʱ�ӣ�10ms=1,000,000��ʱ�����ڣ�
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        key_sync <= 5'b00000;
        key_clean <= 5'b00000;
        key_cnt <= 24'd0;
    end else begin
        // ��һ����ͬ�������źţ���������̬��
        key_sync <= KEY;
        // �ڶ�����������ʱ
        if (key_sync != key_clean) begin
            key_cnt <= 24'd1000000;  // 100MHz * 10ms = 1e6
        end else if (key_cnt > 24'd0) begin
            key_cnt <= key_cnt - 24'd1;
        end else begin
            key_clean <= key_sync;  // ��ʱ����������������İ����ź�
        end
    end
end

// 7. ���뿪�ط����߼���ͬ����������
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        sw_sync <= 8'b00000000;
        sw_clean <= 8'b00000000;
        sw_cnt <= 24'd0;
    end else begin
        // ��һ����ͬ�����뿪���ź�
        sw_sync <= SW;
        // �ڶ�����������ʱ
        if (sw_sync != sw_clean) begin
            sw_cnt <= 24'd1000000;  // 10ms����
        end else if (sw_cnt > 24'd0) begin
            sw_cnt <= sw_cnt - 24'd1;
        end else begin
            sw_clean <= sw_sync;  // ��ʱ���������·�����Ŀ����ź�
        end
    end
end

// 8. ���󵹼�ʱ�߼���100MHzʱ�ӣ�1��=1e8��ʱ�����ڣ�
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        countdown_cnt <= 32'd0;
        countdown_sec <= 4'd10;
        countdown_cfg <= 4'd10;
        countdown_en <= 1'b0;
    end else begin
        // �д�������������ѡ��״̬����������ʱ�����״δ�����
        if (error_type != 3'b000 && current_mode == S_OP_PARAM && !countdown_en) begin
            countdown_en <= 1'b1;
            countdown_cnt <= 32'd100000000 * countdown_cfg;  // 100MHz * N��
            countdown_sec <= countdown_cfg;  // ��ʼʣ������=����ֵ
        end
        // ����ʱ�ڼ䣺�ݼ�������ʵʱ����ʣ������
        if (countdown_en && countdown_cnt > 32'd0) begin
            countdown_cnt <= countdown_cnt - 32'd1;
            countdown_sec <= countdown_cnt / 32'd100000000;  // ʣ������=��ǰ����/1e8
        end
        // ����ʱ����������
        else if (countdown_en && countdown_cnt == 32'd0) begin
            countdown_en <= 1'b0;
            countdown_sec <= countdown_cfg;
            current_mode <= S_OP_PARAM;  // �ص�������ѡ����ʼ�׶�
        end
        // �������Ϸ����˳�����ѡ��״̬�������رյ���ʱ
        if (error_type == 3'b000 || current_mode != S_OP_PARAM) begin
            countdown_en <= 1'b0;
            countdown_sec <= countdown_cfg;
        end
    end
end

// 9. ״̬��ת�߼�������֧��"������ǰģʽ"��
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        current_mode <= S_MENU;
    end else begin
        // ����ʱ�ڼ䣬����������ѡ���������򷵻�
        if (countdown_en) begin
            case (current_mode)
                S_OP_PARAM: begin
                    if (key_clean[0] == 1'b1) begin  // ��S1ȷ����������
                        current_mode <= S_OP_EXEC;
                    end else if (key_clean[2] == 1'b1) begin  // ��S3������������ѡ��
                        current_mode <= S_OP_SELECT;
                        countdown_en <= 1'b0;
                    end else if (key_clean[3] == 1'b1) begin  // ��S4�����˵�
                        current_mode <= S_MENU;
                        countdown_en <= 1'b0;
                    end
                end
                default: current_mode <= current_mode;  // ����״̬����
            endcase
        end else begin
            // �������̣�֧��"������ǰģʽ"��"�������˵�"
            case (current_mode)
                // ���˵���SW5~SW7ѡ��+S1ȷ��
                S_MENU: begin
                    if (key_clean[0] == 1'b1) begin
                        case (sw_clean[7:5])
                            3'b000: current_mode <= S_INPUT;
                            3'b001: current_mode <= S_GEN;
                            3'b010: current_mode <= S_SHOW;
                            3'b011: current_mode <= S_OP_SELECT;
                            default: current_mode <= S_MENU;
                        endcase
                    end else if (key_clean[3] == 1'b1) begin
                        current_mode <= S_MENU;
                    end
                end

                // ����ģʽ��������ɺ�S1/S3�������˵���S2��������
                S_INPUT: begin
                    if (input_done == 1'b1) begin
                        if (key_clean[0] == 1'b1 || key_clean[2] == 1'b1) begin
                            current_mode <= S_MENU;
                        end else if (key_clean[1] == 1'b1) begin  // ������ǰģʽ
                            current_mode <= S_INPUT;
                        end
                    end
                end

                // ����ģʽ��������ģʽ�߼�һ��
                S_GEN: begin
                    if (input_done == 1'b1) begin
                        if (key_clean[0] == 1'b1 || key_clean[2] == 1'b1) begin
                            current_mode <= S_MENU;
                        end else if (key_clean[1] == 1'b1) begin  // ������ǰģʽ
                            current_mode <= S_GEN;
                        end
                    end
                end

                // չʾģʽ��չʾ��ɺ�S1�������˵���S2����չʾ
                S_SHOW: begin
                    if (display_done == 1'b1) begin
                        if (key_clean[0] == 1'b1) begin
                            current_mode <= S_MENU;
                        end else if (key_clean[1] == 1'b1) begin  // ������ǰģʽ
                            current_mode <= S_SHOW;
                        end
                    end
                end

                // ��������ѡ��S1ȷ�ϣ�S3�������˵�
                S_OP_SELECT: begin
                    if (key_clean[0] == 1'b1) begin
                        current_op <= sw_clean[2:0];
                        current_mode <= S_OP_PARAM;
                    end else if (key_clean[2] == 1'b1) begin
                        current_mode <= S_MENU;
                    end
                end

                // ѡ����������S1ȷ�ϣ�S3���أ�S5�л����ѡ��
                S_OP_PARAM: begin
                    if (key_clean[0] == 1'b1) begin
                        if (current_op == OP_SCALAR) begin
                            scalar <= {2'b00, sw_clean[4:3]};  // SW3~SW4ѡ�������0~3��
                        end
                        current_mode <= S_OP_EXEC;
                    end else if (key_clean[2] == 1'b1) begin
                        current_mode <= S_OP_SELECT;
                    end else if (key_clean[4] == 1'b1) begin
                        operand_sel <= 2'b01;  // �л�Ϊϵͳ���ѡ��
                    end
                end

                // ִ�����㣺����Ӧ������ɱ�־
                S_OP_EXEC: begin
                    if (op_done == 1'b1) begin
                        current_mode <= S_RESULT;
                    end
                end

                // չʾ�����S1/S4�����˵���S2������ǰ��������
                S_RESULT: begin
                    if (key_clean[0] == 1'b1 || key_clean[3] == 1'b1) begin
                        current_mode <= S_MENU;
                    end else if (key_clean[1] == 1'b1) begin  // ������ǰ����
                        current_mode <= S_OP_PARAM;
                    end
                end

                S_RETURN: begin
                    current_mode <= S_MENU;
                end

                // �쳣״̬����λ�ؼ��Ĵ����������˵�
                default: begin
                    current_mode <= S_MENU;
                    countdown_en <= 1'b0;
                    operand_sel <= 2'b00;
                    current_op <= OP_TRANS;
                end
            endcase
        end
    end
end

// 10. LED�����߼����ߵ�ƽ������ƥ��Լ���ļ����ţ�
always @(*) begin
    LED = 8'b00000000;  // Ĭ��ȫ��
    case (current_mode)
        S_MENU:      LED[0] = 1'b1;  // LED0=���˵���K3���ţ�
        S_INPUT:     LED[1] = 1'b1;  // LED1=����ģʽ��M1���ţ�
        S_GEN:       LED[2] = 1'b1;  // LED2=����ģʽ��L1���ţ�
        S_SHOW:      LED[3] = 1'b1;  // LED3=չʾģʽ��K6���ţ�
        S_OP_SELECT,
        S_OP_PARAM,
        S_OP_EXEC,
        S_RESULT:    LED[4] = 1'b1;  // LED4=����ģʽ��J5���ţ�
    endcase
    // �д���򵹼�ʱ�ڼ䣬����LED5~LED7��H5��H6��K1���ţ�
    if (error_type != 3'b000 || countdown_en) begin
        LED[5] = 1'b1;
        LED[6] = 1'b1;
        LED[7] = 1'b1;
    end
end

// 11. ����ܿ����߼���16λ��ƥ��Լ���ļ����ţ�
always @(*) begin
    seg_code = {SEG_OFF, SEG_OFF};  // Ĭ��Ϩ��
    if (countdown_en) begin
        // ����ʱ�ڼ䣺��4λ=ʮλ����4λ=��λ
        case (countdown_sec / 4'd10)  // ʮλ��seg_code[15:8]��
            4'd0: seg_code[15:8] = SEG_OFF;
            4'd1: seg_code[15:8] = SEG_1;
            default: seg_code[15:8] = SEG_OFF;
        endcase
        case (countdown_sec % 4'd10)  // ��λ��seg_code[7:0]��
            4'd0: seg_code[7:0] = SEG_0;
            4'd1: seg_code[7:0] = SEG_1;
            4'd2: seg_code[7:0] = SEG_2;
            4'd3: seg_code[7:0] = SEG_3;
            4'd4: seg_code[7:0] = SEG_4;
            4'd5: seg_code[7:0] = SEG_5;
            4'd6: seg_code[7:0] = SEG_6;
            4'd7: seg_code[7:0] = SEG_7;
            4'd8: seg_code[7:0] = SEG_8;
            4'd9: seg_code[7:0] = SEG_9;
            default: seg_code[7:0] = SEG_0;
        endcase
    end else begin
        case (current_mode)
            // ��������ѡ����4λ��ʾ�������ͣ���4λϨ��
            S_OP_SELECT: begin
                case (sw_clean[2:0])
                    OP_TRANS:  seg_code[15:8] = SEG_T;
                    OP_ADD:    seg_code[15:8] = SEG_A;
                    OP_SCALAR: seg_code[15:8] = SEG_B;
                    OP_MUL:    seg_code[15:8] = SEG_C;
                    OP_CONV:   seg_code[15:8] = SEG_J;
                    default:   seg_code[15:8] = SEG_OFF;
                endcase
                seg_code[7:0] = SEG_OFF;
            end
            // ����/����ģʽ����4λ��ʾά�ȣ�SW3~SW4��
            S_INPUT, S_GEN: begin
                case (sw_clean[4:3])
                    2'b00: seg_code[7:0] = SEG_1;  // 1��/��
                    2'b01: seg_code[7:0] = SEG_2;  // 2��/��
                    2'b10: seg_code[7:0] = SEG_3;  // 3��/��
                    2'b11: seg_code[7:0] = SEG_4;  // 4��/��
                    default: seg_code[7:0] = SEG_1;
                endcase
                seg_code[15:8] = SEG_OFF;
            end
            // չʾ�������4λ��ʾ��������4λ��ʾ����
            S_RESULT: begin
                // ������ʾ��result_m=1~5��
                case (result_m)
                    4'd1: seg_code[15:8] = SEG_1;
                    4'd2: seg_code[15:8] = SEG_2;
                    4'd3: seg_code[15:8] = SEG_3;
                    4'd4: seg_code[15:8] = SEG_4;
                    4'd5: seg_code[15:8] = SEG_5;
                    default: seg_code[15:8] = SEG_OFF;
                endcase
                // ������ʾ��result_n=1~5��
                case (result_n)
                    4'd1: seg_code[7:0] = SEG_1;
                    4'd2: seg_code[7:0] = SEG_2;
                    4'd3: seg_code[7:0] = SEG_3;
                    4'd4: seg_code[7:0] = SEG_4;
                    4'd5: seg_code[7:0] = SEG_5;
                    default: seg_code[7:0] = SEG_OFF;
                endcase
            end
        endcase
    end
end

endmodule