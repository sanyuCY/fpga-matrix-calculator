`timescale 1ns / 1ps

module param_config(
    input clk,
    input rst_n,
    input [7:0] uart_rx_data,
    input rx_done,
    output reg [3:0] max_mat_num,    // ÿ�ֹ��������洢����(1~5)
    output reg [7:0] val_min,       // ����Ԫ����Сֵ(-3~20�������ʾ)
    output reg [7:0] val_max,       // ����Ԫ�����ֵ(0~20)
    output reg config_done,         // ������ɱ�־(�ߵ�ƽ����)
    output reg [2:0] error_type     // ��������(000=�޴�,010=ָ���ʽ��,011=�����Ƿ�,100=�洢�����Ƿ�)
);

// ���������������(�����ɶ���)
localparam MIN_NEG3 = 8'd253;  // -3��8λ����
localparam MIN_NEG2 = 8'd254;  // -2��8λ����
localparam MIN_NEG1 = 8'd255;  // -1��8λ����
localparam MAX_VAL  = 8'd20;   // Ԫ�����ֵ����
localparam MIN_VAL  = 8'd0;    // Ԫ��Ĭ����Сֵ

// ָ�����(���洢16�ֽ�ָ��)
reg [7:0] cmd_buf [0:15];
reg [3:0] cmd_cnt;             // ָ���ֽڼ�����
reg cmd_ready;                 // ָ�������ɱ�־

// ��ʱ�Ĵ���(�洢�����еĲ���ֵ)
reg [7:0] new_val_min;
reg [7:0] new_val_max;
reg [3:0] new_max_mat_num;
reg parsing_error;             // ָ����������־

// ״̬����
reg [1:0] state;
localparam IDLE  = 2'b00;      // ����״̬(�ȴ�ָ��)
localparam PARSE = 2'b01;      // ָ�����״̬
localparam CHECK = 2'b10;      // ����У�������״̬

// --- ��integer��������ģ�鼶�������� ---
integer i;
integer comma_idx;  // ����λ������(����rangeָ����)
integer max_len;    // ���ֵ���ֳ���(����rangeָ����)
integer min_idx;    // ��Сֵ��ʼ����(���˿ո���)
// ----------------------------------------

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // ��λ��ʼ�����ָ�Ĭ�ϲ���
        cmd_cnt <= 4'd0;
        cmd_ready <= 1'b0;
        parsing_error <= 1'b0;
        config_done <= 1'b0;
        error_type <= 3'b000;
        state <= IDLE;
        
        // ��ʼ��ָ�����
        for (i = 0; i < 16; i = i + 1) begin
            cmd_buf[i] <= 8'd0;
        end
        
        // ��ʼ����ʱ�Ĵ���(Ĭ�ϲ���)
        new_max_mat_num <= 4'd2;  // Ĭ�ϴ洢2��ͬ������
        new_val_min <= MIN_VAL;   // Ĭ��Ԫ����Сֵ0
        new_val_max <= 8'd9;      // Ĭ��Ԫ�����ֵ9
        
        // ��ʼ������Ĵ���(Ĭ�ϲ���)
        max_mat_num <= 4'd2;
        val_min <= MIN_VAL;
        val_max <= 8'd9;
    end else begin
        case (state)
            // ״̬1������̬������UARTָ��
            IDLE: begin
                config_done <= 1'b0;  // ����������ɱ�־
                error_type <= 3'b000; // �����������
                if (rx_done) begin
                    if (uart_rx_data == 8'h0D) begin  // ��⵽�س���(ָ�����)
                        cmd_ready <= 1'b1;
                        cmd_cnt <= 4'd0;              // ���ü�������׼����һ��ָ��
                        state <= PARSE;
                    end else if (cmd_cnt < 4'd15) begin  // ָ��δ������������������
                        cmd_buf[cmd_cnt] <= uart_rx_data;
                        cmd_cnt <= cmd_cnt + 4'd1;
                    end
                end
            end
            
            // ״̬2������ָ��(x=N �� range=min,max)
            PARSE: begin
                cmd_ready <= 1'b0;
                parsing_error <= 1'b0;
                error_type <= 3'b000;
                
                // ����"x=N"ָ��(����ͬ���������洢����)
                if (cmd_buf[0] == "x" && cmd_buf[1] == "=") begin
                    case (cmd_buf[2])
                        "1": new_max_mat_num <= 4'd1;
                        "2": new_max_mat_num <= 4'd2;
                        "3": new_max_mat_num <= 4'd3;
                        "4": new_max_mat_num <= 4'd4;
                        "5": new_max_mat_num <= 4'd5;
                        default: begin  // �洢��������1~5��Χ
                            parsing_error <= 1'b1;
                            error_type <= 3'b100;
                        end
                    endcase
                end
                // ����"range=min,max"ָ��(����Ԫ��ֵ��Χ)
                else if (cmd_buf[0] == "r" && cmd_buf[1] == "a" && 
                         cmd_buf[2] == "n" && cmd_buf[3] == "g" && 
                         cmd_buf[4] == "e" && cmd_buf[5] == "=") begin
                    // ����1���ҵ����ŷָ���
                    comma_idx = 6;
                    while (comma_idx < 15 && cmd_buf[comma_idx] != ",") begin
                        comma_idx = comma_idx + 1;
                    end
                    
                    if (comma_idx >= 15) begin  // δ�ҵ����ţ�ָ���ʽ����
                        parsing_error <= 1'b1;
                        error_type <= 3'b010;
                    end else begin
                        // ����2��������Сֵ(���˿ո�֧�ָ���)
                        min_idx = 6;
                        while (min_idx < comma_idx && cmd_buf[min_idx] == " ") begin  // �����ո�
                            min_idx = min_idx + 1;
                        end
                        
                        if (cmd_buf[min_idx] == "-") begin  // ������(-1~-3)
                            case (cmd_buf[min_idx+1])
                                "1": new_val_min <= MIN_NEG1;
                                "2": new_val_min <= MIN_NEG2;
                                "3": new_val_min <= MIN_NEG3;
                                default: begin  // ��������-3��Χ
                                    parsing_error <= 1'b1;
                                    error_type <= 3'b011;
                                end
                            endcase
                        end else begin  // ��������(0~20)
                            if (comma_idx - min_idx == 1) begin  // 1λ����(��"5,")
                                new_val_min <= cmd_buf[min_idx] - 8'h30;
                            end else if (comma_idx - min_idx == 2) begin  // 2λ����(��"15,")
                                new_val_min <= (cmd_buf[min_idx] - 8'h30) * 10 + (cmd_buf[min_idx+1] - 8'h30);
                            end else begin  // ����λ������
                                parsing_error <= 1'b1;
                                error_type <= 3'b011;
                            end
                        end
                        
                        // ����3���������ֵ(���ź󣬽�֧������0~20)
                        max_len = cmd_cnt - comma_idx - 1;  // ���ֵ���ֳ���
                        if (max_len == 1) begin  // 1λ���ֵ(��",5")
                            new_val_max <= cmd_buf[comma_idx+1] - 8'h30;
                        end else if (max_len == 2) begin  // 2λ���ֵ(��",15")
                            new_val_max <= (cmd_buf[comma_idx+1] - 8'h30) * 10 + (cmd_buf[comma_idx+2] - 8'h30);
                        end else begin  // ���ֵλ������
                            parsing_error <= 1'b1;
                            error_type <= 3'b011;
                        end
                    end
                end
                // δָ֪���ʽ
                else begin
                    parsing_error <= 1'b1;
                    error_type <= 3'b010;
                end
                
                state <= CHECK;  // �������У��״̬
            end
            
            // ״̬3�������Ϸ���У�������
            CHECK: begin
                if (!parsing_error) begin
                    // �Ӳ���1�����²���(����ָ������)
                    if (cmd_buf[0] == "x") begin  // ����x=Nָ��
                        max_mat_num <= new_max_mat_num;
                        // ����У��洢����(ȷ��1~5)
                        if (max_mat_num < 4'd1) begin
                            max_mat_num <= 4'd1;
                            error_type <= 3'b100;
                        end else if (max_mat_num > 4'd5) begin
                            max_mat_num <= 4'd5;
                            error_type <= 3'b100;
                        end
                    end else if (cmd_buf[0] == "r") begin  // ����rangeָ��
                        val_min <= new_val_min;
                        val_max <= new_val_max;
                        // ����У��Ԫ�ط�Χ
                        // У��val_min��-3(253)~20
                        if (val_min < MIN_NEG3 || val_min > MAX_VAL) begin
                            val_min <= MIN_VAL;
                            error_type <= 3'b011;
                        end
                        // У��val_max��0~20
                        if (val_max < MIN_VAL || val_max > MAX_VAL) begin
                            val_max <= 8'd9;
                            error_type <= 3'b011;
                        end
                        // У��val_max >= val_min(����ָ�Ĭ��0~9)
                        if (val_max < val_min) begin
                            val_min <= MIN_VAL;
                            val_max <= 8'd9;
                            error_type <= 3'b011;
                        end
                    end
                    
                    // �Ӳ���2������������ɱ�־(�޴���ʱ)
                    if (error_type == 3'b000) begin
                        config_done <= 1'b1;
                    end
                end
                
                // �Ӳ���3��������������ʱ�Ĵ���
                cmd_cnt <= 4'd0;
                for (i = 0; i < 16; i = i + 1) begin
                    cmd_buf[i] <= 8'd0;
                end
                new_val_min <= MIN_VAL;   // ������ʱ��Сֵ
                new_val_max <= 8'd9;      // ������ʱ���ֵ
                new_max_mat_num <= 4'd2;  // ������ʱ�洢����
                
                state <= IDLE;  // ���ؿ���̬���ȴ���һ��ָ��
            end
        endcase
    end
end

endmodule


