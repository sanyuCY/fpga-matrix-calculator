//�����������ģ��
// ģ�鹦�ܣ�����UART��������ľ������ݣ����ά��/Ԫ�غϷ��Լ�⣬����ṹ����������
module matrix_input(
    input clk,
    input rst_n,// �͵�ƽ��λ��0=��λ��1=����������
    //����UARTģ��
    input [7:0] uart_rx_data, // UART���յĵ��ֽ����ݣ�ASCII�룬8λ��
    input rx_done,      // UART���ֽڽ�����ɱ�־���ߵ�ƽ��Ч������1��ʱ�ӣ�
    // ����FSMģ��
    input [3:0] val_min,
    input [3:0]  val_max,
    //�����λ�Ա㸲�ǵ�15
    // ������洢/����ģ��ľ�������
    output reg [3:0] mat_m,
    output reg [3:0] mat_n, // ���ڶԽ�
    output reg [3:0] mat_data [0:4][0:4], // 5��5��ά����
    // �����FSMģ���״̬or�����־
    output reg input_done, // ���������ɱ�־���ߵ�ƽ��Ч������1��ʱ�ӣ�
    output reg [2:0] error_type  // �������ͣ�3λ���ͽӿ��ֲ�һ�£�000=�޴�001=ά�ȴ�011=Ԫ��ֵ��
);
// 1. ״̬�����壨����״̬��FSM�����ƽ������̣�
// localprarm��ߴ���ɶ���ͬʱ����ά���ɱ�
localparam S_WAIT = 3'b000; // �ȴ�UART��������
localparam S_PARSE_M = 3'b001; // ������������m
localparam S_PARSE_N = 3'b010; // ������������n
localparam S_PARSE_DATA= 3'b011; // ��������Ԫ��
localparam S_CHECK = 3'b100; // �Ϸ��Լ��
localparam S_DONE = 3'b101; // ������ɣ�������
// 2. ״̬���Ĵ������洢��ǰ״̬��
reg [2:0] curr_state;  // ��ǰ״̬
reg [2:0] next_state;  // ��һ״̬������ʽ״̬��������ȶ��ԣ�
// 3. ��ʱ�洢�Ĵ���������ֱ�Ӹ�������Ĵ�����
reg [3:0] m_temp;      // ������ʱ���棨������ɺ��ٸ�ֵ��mat_m��
reg [3:0] n_temp;      // ������ʱ����
reg [3:0] data_temp [0:4][0:4]; // Ԫ����ʱ���棨��������������Ч���ݣ�
// 4. �����Ĵ�����ͳ���ѽ�����Ԫ�ظ�����
reg [4:0]  data_cnt;    // Ԫ�ؼ�������0~24��5��5=25��Ԫ�أ�
// ���ܣ���ʱ�������ظ��µ�ǰ״̬����λʱ�ص��ȴ�״̬��
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        curr_state <= S_WAIT; // ��λ���ʼ״̬���ȴ�
    end else begin
        curr_state <= next_state; // �Ǹ�λʱ������Ϊ��һ״̬
    end
end
// ���ܣ����ݵ�ǰ״̬+����������������һ״̬����ʱ�򣬴��߼��жϣ�
always @(*) begin
    next_state = curr_state; // Ĭ�ϱ��ֵ�ǰ״̬���������������ɣ�
    case(curr_state)
        S_WAIT: begin
            // ����������UART�յ���һ���ֽڣ�����m��
            if(rx_done) begin
                next_state = S_PARSE_M;
            end
        end
        S_PARSE_M: begin
            // ����������UART�յ��ڶ����ֽڣ�����n��
            if(rx_done) begin
                next_state = S_PARSE_N;
            end
        end
        S_PARSE_N: begin
            // ����������UART�յ��������ֽڣ���һ��Ԫ�أ�
            if(rx_done) begin
                next_state = S_PARSE_DATA;
            end
        end
        S_PARSE_DATA: begin
            // ����������Ԫ�ؽ�����ɣ��������ﵽm��n-1�����յ����һ��Ԫ��
            if(rx_done && (data_cnt == m_temp * n_temp - 1)) begin
                next_state = S_CHECK;
            end
        end
        S_CHECK: begin
            // �Ϸ��Լ����ɺ�ֱ�ӽ������״̬
            next_state = S_DONE;
        end
        S_DONE: begin
            // ��ɺ�ص��ȴ�״̬��׼����һ�ν���
            next_state = S_WAIT;
        end
        default: begin
            next_state = S_WAIT; // �쳣״̬�ص��ȴ������³����
        end
    endcase
end
// ���ܣ��ڲ�ͬ״̬�£�����UART���ݵ���ʱ�Ĵ���
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        // ��λ�����������ʱ�Ĵ����ͼ�����
        m_temp <= 4'd0;
        n_temp <= 4'd0;
        data_temp[0][0] <= 4'd0;
        data_temp[0][1] <= 4'd0;
        data_temp[0][2] <= 4'd0;
        data_temp[0][3] <= 4'd0;
        data_temp[0][4] <= 4'd0;
        data_temp[1][0] <= 4'd0;
        data_temp[1][1] <= 4'd0;
        data_temp[1][2] <= 4'd0;
        data_temp[1][3] <= 4'd0;
        data_temp[1][4] <= 4'd0;
        data_temp[2][0] <= 4'd0;
        data_temp[2][1] <= 4'd0;
        data_temp[2][2] <= 4'd0;
        data_temp[2][3] <= 4'd0;
        data_temp[2][4] <= 4'd0;
        data_temp[3][0] <= 4'd0;
        data_temp[3][1] <= 4'd0;
        data_temp[3][2] <= 4'd0;
        data_temp[3][3] <= 4'd0;
        data_temp[3][4] <= 4'd0;
        data_temp[4][0] <= 4'd0;
        data_temp[4][1] <= 4'd0;
        data_temp[4][2] <= 4'd0;
        data_temp[4][3] <= 4'd0;
        data_temp[4][4] <= 4'd0;
        data_cnt <= 5'd0;
    end else begin
        case(curr_state)
            S_PARSE_M: begin
                // ASCII0-9���������λΪ���ֱ���
                if(rx_done) begin
                    m_temp <= uart_rx_data[3:0]; // 8'h32�ĵ�4λ��2�����ASCII������ת��
                end
            end
            S_PARSE_N: begin
                // ��������n���������߼�һ��
                if(rx_done) begin
                    n_temp <= uart_rx_data[3:0];
                end
            end
            S_PARSE_DATA: begin
                // ����Ԫ�أ������������洢����ʱ����
                if(rx_done) begin
                    // Ԫ���������ҵ��ڼ��еڼ���
                    data_temp[data_cnt / n_temp][data_cnt % n_temp] <= uart_rx_data[3:0];
                    data_cnt <= data_cnt + 1'b1; // ����������
                end
            end
            S_DONE: begin
                // ������ɺ����ü�����
                data_cnt <= 5'd0;
            end
            default: begin
                // ����״̬������ʱ�Ĵ�������
                m_temp <= m_temp;
                n_temp <= n_temp;
                data_cnt <= data_cnt;
            end
        endcase
    end
end
integer i, j;
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        // ��λ���������Ĵ����ͱ�־
        mat_m <= 4'd0;
        mat_n <= 4'd0;
        mat_data[0][0] <= 4'd0;
        mat_data[0][1] <= 4'd0;
        mat_data[0][2] <= 4'd0;
        mat_data[0][3] <= 4'd0;
        mat_data[0][4] <= 4'd0;
        mat_data[1][0] <= 4'd0;
        mat_data[1][1] <= 4'd0;
        mat_data[1][2] <= 4'd0;
        mat_data[1][3] <= 4'd0;
        mat_data[1][4] <= 4'd0;
        mat_data[2][0] <= 4'd0;
        mat_data[2][1] <= 4'd0;
        mat_data[2][2] <= 4'd0;
        mat_data[2][3] <= 4'd0;
        mat_data[2][4] <= 4'd0;
        mat_data[3][0] <= 4'd0;
        mat_data[3][1] <= 4'd0;
        mat_data[3][2] <= 4'd0;
        mat_data[3][3] <= 4'd0;
        mat_data[3][4] <= 4'd0;
        mat_data[4][0] <= 4'd0;
        mat_data[4][1] <= 4'd0;
        mat_data[4][2] <= 4'd0;
        mat_data[4][3] <= 4'd0;
        mat_data[4][4] <= 4'd0;
        input_done <= 1'b0;
        error_type <= 3'b000;
    end else begin
        case(curr_state)
            S_CHECK: begin
                // ��ʼ����������Ϊ�޴�
                error_type <= 3'b000;
                
                // ���ά�ȺϷ��ԣ�1~5��
                if(m_temp < 4'd1 || m_temp > 4'd5 || n_temp < 4'd1 || n_temp > 4'd5) begin
                    error_type <= 3'b001; // ά�ȴ���001
                end else begin
                    // �ڶ��������Ԫ��ֵ�Ϸ��ԣ�val_min~val_max��
                    for(i=0; i<m_temp; i=i+1) begin 
                        for(j=0; j<n_temp; j=j+1) begin 
                            if(data_temp[i][j] < val_min || data_temp[i][j] > val_max) begin
                                error_type <= 3'b011; // Ԫ��ֵ����011
                            end
                        end
                    end
                end
            end
            S_DONE: begin
                // �޴���ʱ������ʱ���ݸ�ֵ������Ĵ���
                if(error_type == 3'b000) begin
                    mat_m <= m_temp;
                    mat_n <= n_temp;
                    for(i=0; i<m_temp; i=i+1) begin
                        for(j=0; j<n_temp; j=j+1) begin
                            mat_data[i][j] <= data_temp[i][j];
                        end
                    end
                end else begin
                    // �д���ʱ������������������Ƿ����ݣ�
                    mat_m <= 4'd0;
                    mat_n <= 4'd0;
                    mat_data[0][0] <= 4'd0;
                    mat_data[0][1] <= 4'd0;
                    mat_data[0][2] <= 4'd0;
                    mat_data[0][3] <= 4'd0;
                    mat_data[0][4] <= 4'd0;
                    mat_data[1][0] <= 4'd0;
                    mat_data[1][1] <= 4'd0;
                    mat_data[1][2] <= 4'd0;
                    mat_data[1][3] <= 4'd0;
                    mat_data[1][4] <= 4'd0;
                    mat_data[2][0] <= 4'd0;
                    mat_data[2][1] <= 4'd0;
                    mat_data[2][2] <= 4'd0;
                    mat_data[2][3] <= 4'd0;
                    mat_data[2][4] <= 4'd0;
                    mat_data[3][0] <= 4'd0;
                    mat_data[3][1] <= 4'd0;
                    mat_data[3][2] <= 4'd0;
                    mat_data[3][3] <= 4'd0;
                    mat_data[3][4] <= 4'd0;
                    mat_data[4][0] <= 4'd0;
                    mat_data[4][1] <= 4'd0;
                    mat_data[4][2] <= 4'd0;
                    mat_data[4][3] <= 4'd0;
                    mat_data[4][4] <= 4'd0;
                end
                // ��λ��ɱ�־������FSMģ�������ɣ�
                input_done <= 1'b1;
            end
            default: begin
                // ����״̬�������ɱ�־�����ִ�������
                input_done <= 1'b0;
                error_type <= error_type;
            end
        endcase
    end
end
endmodule