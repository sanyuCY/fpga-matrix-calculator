`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////
// Module: matrix_storage - �����棨Vivado 2017���ݣ�
// ���ܣ�
//   1. ��������(m*n)����洢
//   2. ÿ�ֹ�����洢 max_mat_num ������
//   3. ͬ�����󳬳�����ʱ��������ɵģ���ת���ǣ�
//   4. spec_count_flat ���ÿ�ֹ��ľ�������ͳ��
//////////////////////////////////////////////////////////////////////////////

module matrix_storage (
    input wire clk,
    input wire rst_n,
    input wire [3:0] max_mat_num,           // ÿ�ֹ�����洢�ľ�������Ĭ��2��
    
    // ����ģ��ӿ�
    input wire [3:0] input_mat_m,
    input wire [3:0] input_mat_n,
    input wire [199:0] input_mat_data,
    input wire input_store_en,
    
    // ����ģ��ӿ�
    input wire [3:0] gen_mat_m,
    input wire [3:0] gen_mat_n,
    input wire [199:0] gen_mat_data,
    input wire gen_store_en,
    
    // ��ȡ�ӿ�
    input wire [3:0] read_idx,
    input wire read_en,
    
    // ��������д洢�����չƽ����
    output wire [39:0] stored_mat_m_flat,
    output wire [39:0] stored_mat_n_flat,
    output wire [39:0] stored_mat_id_flat,
    output wire [1999:0] stored_mat_flat,
    output reg [3:0] total_mat_count,
    
    // ��ȡ���
    output reg [3:0] read_out_m,
    output reg [3:0] read_out_n,
    output reg [199:0] read_out_data,
    output reg [3:0] read_out_id,
    output reg read_valid,
    output reg read_done,
    
    // ���ͳ�ƣ�25�ֹ��(1-5 * 1-5)��ÿ��4bit����
    output wire [99:0] spec_count_flat,
    
    output reg [2:0] error_type
);

    //==========================================================================
    // �洢�ṹ��10�������λ��ʹ�ö����Ĵ�����Vivado 2017���ݣ�
    //==========================================================================
    reg [3:0] mat_m_0, mat_m_1, mat_m_2, mat_m_3, mat_m_4;
    reg [3:0] mat_m_5, mat_m_6, mat_m_7, mat_m_8, mat_m_9;
    reg [3:0] mat_n_0, mat_n_1, mat_n_2, mat_n_3, mat_n_4;
    reg [3:0] mat_n_5, mat_n_6, mat_n_7, mat_n_8, mat_n_9;
    reg [3:0] mat_id_0, mat_id_1, mat_id_2, mat_id_3, mat_id_4;
    reg [3:0] mat_id_5, mat_id_6, mat_id_7, mat_id_8, mat_id_9;
    reg [199:0] mat_data_0, mat_data_1, mat_data_2, mat_data_3, mat_data_4;
    reg [199:0] mat_data_5, mat_data_6, mat_data_7, mat_data_8, mat_data_9;
    reg mat_valid_0, mat_valid_1, mat_valid_2, mat_valid_3, mat_valid_4;
    reg mat_valid_5, mat_valid_6, mat_valid_7, mat_valid_8, mat_valid_9;
    
    reg [3:0] next_id;
    
    //==========================================================================
    // ÿ�ֹ��(m,n)�ļ�����
    // ������� = (m-1)*5 + (n-1)����Χ0-24
    //==========================================================================
    reg [3:0] spec_count_0,  spec_count_1,  spec_count_2,  spec_count_3,  spec_count_4;
    reg [3:0] spec_count_5,  spec_count_6,  spec_count_7,  spec_count_8,  spec_count_9;
    reg [3:0] spec_count_10, spec_count_11, spec_count_12, spec_count_13, spec_count_14;
    reg [3:0] spec_count_15, spec_count_16, spec_count_17, spec_count_18, spec_count_19;
    reg [3:0] spec_count_20, spec_count_21, spec_count_22, spec_count_23, spec_count_24;
    
    //==========================================================================
    // ���չƽ������ԭ�ӿڣ�
    //==========================================================================
    assign stored_mat_m_flat = {mat_m_9, mat_m_8, mat_m_7, mat_m_6, mat_m_5,
                                mat_m_4, mat_m_3, mat_m_2, mat_m_1, mat_m_0};
    assign stored_mat_n_flat = {mat_n_9, mat_n_8, mat_n_7, mat_n_6, mat_n_5,
                                mat_n_4, mat_n_3, mat_n_2, mat_n_1, mat_n_0};
    assign stored_mat_id_flat = {mat_id_9, mat_id_8, mat_id_7, mat_id_6, mat_id_5,
                                 mat_id_4, mat_id_3, mat_id_2, mat_id_1, mat_id_0};
    assign stored_mat_flat = {mat_data_9, mat_data_8, mat_data_7, mat_data_6, mat_data_5,
                              mat_data_4, mat_data_3, mat_data_2, mat_data_1, mat_data_0};
    
    // ������չƽ���
    assign spec_count_flat = {spec_count_24, spec_count_23, spec_count_22, spec_count_21, spec_count_20,
                              spec_count_19, spec_count_18, spec_count_17, spec_count_16, spec_count_15,
                              spec_count_14, spec_count_13, spec_count_12, spec_count_11, spec_count_10,
                              spec_count_9,  spec_count_8,  spec_count_7,  spec_count_6,  spec_count_5,
                              spec_count_4,  spec_count_3,  spec_count_2,  spec_count_1,  spec_count_0};
    
    //==========================================================================
    // �ڲ��ź�
    //==========================================================================
    wire store_en;
    wire [3:0] store_m, store_n;
    wire [199:0] store_data;
    wire [4:0] spec_idx;                    // ������� = (m-1)*5 + (n-1)
    
    assign store_en = input_store_en | gen_store_en;
    assign store_m = input_store_en ? input_mat_m : gen_mat_m;
    assign store_n = input_store_en ? input_mat_n : gen_mat_n;
    assign store_data = input_store_en ? input_mat_data : gen_mat_data;
    assign spec_idx = (store_m - 1) * 5 + (store_n - 1);
    
    //==========================================================================
    // ����ͬ���������������ɲ�λ
    //==========================================================================
    reg [3:0] match_count;
    reg [3:0] oldest_slot;
    reg [3:0] oldest_id;
    reg [3:0] empty_slot;
    reg found_empty;
    reg [3:0] target_slot;
    reg need_overwrite;
    reg [4:0] old_spec_idx;                 // �����ǲ�λ��ԭ�������
    
    // ��ʱ�������ڱ���
    wire match_0, match_1, match_2, match_3, match_4;
    wire match_5, match_6, match_7, match_8, match_9;
    
    assign match_0 = mat_valid_0 && (mat_m_0 == store_m) && (mat_n_0 == store_n);
    assign match_1 = mat_valid_1 && (mat_m_1 == store_m) && (mat_n_1 == store_n);
    assign match_2 = mat_valid_2 && (mat_m_2 == store_m) && (mat_n_2 == store_n);
    assign match_3 = mat_valid_3 && (mat_m_3 == store_m) && (mat_n_3 == store_n);
    assign match_4 = mat_valid_4 && (mat_m_4 == store_m) && (mat_n_4 == store_n);
    assign match_5 = mat_valid_5 && (mat_m_5 == store_m) && (mat_n_5 == store_n);
    assign match_6 = mat_valid_6 && (mat_m_6 == store_m) && (mat_n_6 == store_n);
    assign match_7 = mat_valid_7 && (mat_m_7 == store_m) && (mat_n_7 == store_n);
    assign match_8 = mat_valid_8 && (mat_m_8 == store_m) && (mat_n_8 == store_n);
    assign match_9 = mat_valid_9 && (mat_m_9 == store_m) && (mat_n_9 == store_n);
    
    // ����߼�������Ŀ���λ
    always @(*) begin
        // ����ƥ������
        match_count = {3'd0, match_0} + {3'd0, match_1} + {3'd0, match_2} + 
                      {3'd0, match_3} + {3'd0, match_4} + {3'd0, match_5} + 
                      {3'd0, match_6} + {3'd0, match_7} + {3'd0, match_8} + {3'd0, match_9};
        
        // ���ҿղ�λ������ѡ������С�ģ�
        found_empty = 1'b0;
        empty_slot = 4'd0;
        if (!mat_valid_0) begin found_empty = 1'b1; empty_slot = 4'd0; end
        else if (!mat_valid_1) begin found_empty = 1'b1; empty_slot = 4'd1; end
        else if (!mat_valid_2) begin found_empty = 1'b1; empty_slot = 4'd2; end
        else if (!mat_valid_3) begin found_empty = 1'b1; empty_slot = 4'd3; end
        else if (!mat_valid_4) begin found_empty = 1'b1; empty_slot = 4'd4; end
        else if (!mat_valid_5) begin found_empty = 1'b1; empty_slot = 4'd5; end
        else if (!mat_valid_6) begin found_empty = 1'b1; empty_slot = 4'd6; end
        else if (!mat_valid_7) begin found_empty = 1'b1; empty_slot = 4'd7; end
        else if (!mat_valid_8) begin found_empty = 1'b1; empty_slot = 4'd8; end
        else if (!mat_valid_9) begin found_empty = 1'b1; empty_slot = 4'd9; end
        
        // ����ͬ�����ID��С����ɣ��Ĳ�λ
        oldest_slot = 4'd0;
        oldest_id = 4'd15;
        
        if (match_0 && mat_id_0 < oldest_id) begin oldest_id = mat_id_0; oldest_slot = 4'd0; end
        if (match_1 && mat_id_1 < oldest_id) begin oldest_id = mat_id_1; oldest_slot = 4'd1; end
        if (match_2 && mat_id_2 < oldest_id) begin oldest_id = mat_id_2; oldest_slot = 4'd2; end
        if (match_3 && mat_id_3 < oldest_id) begin oldest_id = mat_id_3; oldest_slot = 4'd3; end
        if (match_4 && mat_id_4 < oldest_id) begin oldest_id = mat_id_4; oldest_slot = 4'd4; end
        if (match_5 && mat_id_5 < oldest_id) begin oldest_id = mat_id_5; oldest_slot = 4'd5; end
        if (match_6 && mat_id_6 < oldest_id) begin oldest_id = mat_id_6; oldest_slot = 4'd6; end
        if (match_7 && mat_id_7 < oldest_id) begin oldest_id = mat_id_7; oldest_slot = 4'd7; end
        if (match_8 && mat_id_8 < oldest_id) begin oldest_id = mat_id_8; oldest_slot = 4'd8; end
        if (match_9 && mat_id_9 < oldest_id) begin oldest_id = mat_id_9; oldest_slot = 4'd9; end
        
        // ����Ŀ���λ
        if (match_count >= max_mat_num && match_count > 4'd0) begin
            // ͬ����Ѵ����ޣ���Ҫ������ɵ�ͬ������
            need_overwrite = 1'b1;
            target_slot = oldest_slot;
        end
        else if (found_empty) begin
            // �пղ�λ��ʹ�ÿղ�λ��������
            need_overwrite = 1'b0;
            target_slot = empty_slot;
        end
        else if (match_count > 4'd0) begin
            // û�пղ�λ�����ù���о��󣨼�ʹδ�����ޣ�
            // ���ȸ���ͬ�����ɵľ���
            need_overwrite = 1'b1;
            target_slot = oldest_slot;
        end
        else begin
            // û�пղ�λ���Ҹù��û���κξ���
            // ��Ҫ�����������ľ������ڳ��ռ䣨ȫ����ɣ�
            need_overwrite = 1'b0;  // ��������������������spec_count��
            target_slot = 4'd0;
            oldest_id = 4'd15;
            
            // ��ȫ����ɵĲ�λ
            if (mat_valid_0 && mat_id_0 < oldest_id) begin oldest_id = mat_id_0; target_slot = 4'd0; end
            if (mat_valid_1 && mat_id_1 < oldest_id) begin oldest_id = mat_id_1; target_slot = 4'd1; end
            if (mat_valid_2 && mat_id_2 < oldest_id) begin oldest_id = mat_id_2; target_slot = 4'd2; end
            if (mat_valid_3 && mat_id_3 < oldest_id) begin oldest_id = mat_id_3; target_slot = 4'd3; end
            if (mat_valid_4 && mat_id_4 < oldest_id) begin oldest_id = mat_id_4; target_slot = 4'd4; end
            if (mat_valid_5 && mat_id_5 < oldest_id) begin oldest_id = mat_id_5; target_slot = 4'd5; end
            if (mat_valid_6 && mat_id_6 < oldest_id) begin oldest_id = mat_id_6; target_slot = 4'd6; end
            if (mat_valid_7 && mat_id_7 < oldest_id) begin oldest_id = mat_id_7; target_slot = 4'd7; end
            if (mat_valid_8 && mat_id_8 < oldest_id) begin oldest_id = mat_id_8; target_slot = 4'd8; end
            if (mat_valid_9 && mat_id_9 < oldest_id) begin oldest_id = mat_id_9; target_slot = 4'd9; end
        end
        
        // ���㱻���ǲ�λ��ԭ�������
        case (target_slot)
            4'd0: old_spec_idx = (mat_m_0 - 1) * 5 + (mat_n_0 - 1);
            4'd1: old_spec_idx = (mat_m_1 - 1) * 5 + (mat_n_1 - 1);
            4'd2: old_spec_idx = (mat_m_2 - 1) * 5 + (mat_n_2 - 1);
            4'd3: old_spec_idx = (mat_m_3 - 1) * 5 + (mat_n_3 - 1);
            4'd4: old_spec_idx = (mat_m_4 - 1) * 5 + (mat_n_4 - 1);
            4'd5: old_spec_idx = (mat_m_5 - 1) * 5 + (mat_n_5 - 1);
            4'd6: old_spec_idx = (mat_m_6 - 1) * 5 + (mat_n_6 - 1);
            4'd7: old_spec_idx = (mat_m_7 - 1) * 5 + (mat_n_7 - 1);
            4'd8: old_spec_idx = (mat_m_8 - 1) * 5 + (mat_n_8 - 1);
            4'd9: old_spec_idx = (mat_m_9 - 1) * 5 + (mat_n_9 - 1);
            default: old_spec_idx = 5'd0;
        endcase
    end
    
    //==========================================================================
    // ���洢�߼�
    //==========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // ��λ���д洢
            next_id <= 4'd1;
            total_mat_count <= 4'd0;
            error_type <= 3'd0;
            read_valid <= 1'b0;
            read_done <= 1'b0;
            read_out_m <= 4'd0;
            read_out_n <= 4'd0;
            read_out_id <= 4'd0;
            read_out_data <= 200'd0;
            
            // �����λ��λ
            mat_m_0 <= 4'd0; mat_m_1 <= 4'd0; mat_m_2 <= 4'd0; mat_m_3 <= 4'd0; mat_m_4 <= 4'd0;
            mat_m_5 <= 4'd0; mat_m_6 <= 4'd0; mat_m_7 <= 4'd0; mat_m_8 <= 4'd0; mat_m_9 <= 4'd0;
            mat_n_0 <= 4'd0; mat_n_1 <= 4'd0; mat_n_2 <= 4'd0; mat_n_3 <= 4'd0; mat_n_4 <= 4'd0;
            mat_n_5 <= 4'd0; mat_n_6 <= 4'd0; mat_n_7 <= 4'd0; mat_n_8 <= 4'd0; mat_n_9 <= 4'd0;
            mat_id_0 <= 4'd0; mat_id_1 <= 4'd0; mat_id_2 <= 4'd0; mat_id_3 <= 4'd0; mat_id_4 <= 4'd0;
            mat_id_5 <= 4'd0; mat_id_6 <= 4'd0; mat_id_7 <= 4'd0; mat_id_8 <= 4'd0; mat_id_9 <= 4'd0;
            mat_data_0 <= 200'd0; mat_data_1 <= 200'd0; mat_data_2 <= 200'd0;
            mat_data_3 <= 200'd0; mat_data_4 <= 200'd0; mat_data_5 <= 200'd0;
            mat_data_6 <= 200'd0; mat_data_7 <= 200'd0; mat_data_8 <= 200'd0; mat_data_9 <= 200'd0;
            mat_valid_0 <= 1'b0; mat_valid_1 <= 1'b0; mat_valid_2 <= 1'b0;
            mat_valid_3 <= 1'b0; mat_valid_4 <= 1'b0; mat_valid_5 <= 1'b0;
            mat_valid_6 <= 1'b0; mat_valid_7 <= 1'b0; mat_valid_8 <= 1'b0; mat_valid_9 <= 1'b0;
            
            // ��������λ
            spec_count_0  <= 4'd0; spec_count_1  <= 4'd0; spec_count_2  <= 4'd0;
            spec_count_3  <= 4'd0; spec_count_4  <= 4'd0; spec_count_5  <= 4'd0;
            spec_count_6  <= 4'd0; spec_count_7  <= 4'd0; spec_count_8  <= 4'd0;
            spec_count_9  <= 4'd0; spec_count_10 <= 4'd0; spec_count_11 <= 4'd0;
            spec_count_12 <= 4'd0; spec_count_13 <= 4'd0; spec_count_14 <= 4'd0;
            spec_count_15 <= 4'd0; spec_count_16 <= 4'd0; spec_count_17 <= 4'd0;
            spec_count_18 <= 4'd0; spec_count_19 <= 4'd0; spec_count_20 <= 4'd0;
            spec_count_21 <= 4'd0; spec_count_22 <= 4'd0; spec_count_23 <= 4'd0;
            spec_count_24 <= 4'd0;
        end
        else begin
            read_done <= 1'b0;
            error_type <= 3'd0;
            
            //==================================================================
            // �洢������
            //==================================================================
            if (store_en) begin
                // д��Ŀ���λ
                case (target_slot)
                    4'd0: begin
                        mat_m_0 <= store_m; mat_n_0 <= store_n;
                        mat_data_0 <= store_data; mat_id_0 <= next_id;
                        mat_valid_0 <= 1'b1;
                    end
                    4'd1: begin
                        mat_m_1 <= store_m; mat_n_1 <= store_n;
                        mat_data_1 <= store_data; mat_id_1 <= next_id;
                        mat_valid_1 <= 1'b1;
                    end
                    4'd2: begin
                        mat_m_2 <= store_m; mat_n_2 <= store_n;
                        mat_data_2 <= store_data; mat_id_2 <= next_id;
                        mat_valid_2 <= 1'b1;
                    end
                    4'd3: begin
                        mat_m_3 <= store_m; mat_n_3 <= store_n;
                        mat_data_3 <= store_data; mat_id_3 <= next_id;
                        mat_valid_3 <= 1'b1;
                    end
                    4'd4: begin
                        mat_m_4 <= store_m; mat_n_4 <= store_n;
                        mat_data_4 <= store_data; mat_id_4 <= next_id;
                        mat_valid_4 <= 1'b1;
                    end
                    4'd5: begin
                        mat_m_5 <= store_m; mat_n_5 <= store_n;
                        mat_data_5 <= store_data; mat_id_5 <= next_id;
                        mat_valid_5 <= 1'b1;
                    end
                    4'd6: begin
                        mat_m_6 <= store_m; mat_n_6 <= store_n;
                        mat_data_6 <= store_data; mat_id_6 <= next_id;
                        mat_valid_6 <= 1'b1;
                    end
                    4'd7: begin
                        mat_m_7 <= store_m; mat_n_7 <= store_n;
                        mat_data_7 <= store_data; mat_id_7 <= next_id;
                        mat_valid_7 <= 1'b1;
                    end
                    4'd8: begin
                        mat_m_8 <= store_m; mat_n_8 <= store_n;
                        mat_data_8 <= store_data; mat_id_8 <= next_id;
                        mat_valid_8 <= 1'b1;
                    end
                    4'd9: begin
                        mat_m_9 <= store_m; mat_n_9 <= store_n;
                        mat_data_9 <= store_data; mat_id_9 <= next_id;
                        mat_valid_9 <= 1'b1;
                    end
                    default: ;
                endcase
                
                // ����ID
                next_id <= next_id + 4'd1;
                
                // ���������͹�����
                if (!need_overwrite && found_empty) begin
                    // ���1��ʹ�ÿղ�λ����������+1���¹�����+1
                    total_mat_count <= total_mat_count + 4'd1;
                    
                    case (spec_idx)
                        5'd0:  spec_count_0  <= spec_count_0  + 4'd1;
                        5'd1:  spec_count_1  <= spec_count_1  + 4'd1;
                        5'd2:  spec_count_2  <= spec_count_2  + 4'd1;
                        5'd3:  spec_count_3  <= spec_count_3  + 4'd1;
                        5'd4:  spec_count_4  <= spec_count_4  + 4'd1;
                        5'd5:  spec_count_5  <= spec_count_5  + 4'd1;
                        5'd6:  spec_count_6  <= spec_count_6  + 4'd1;
                        5'd7:  spec_count_7  <= spec_count_7  + 4'd1;
                        5'd8:  spec_count_8  <= spec_count_8  + 4'd1;
                        5'd9:  spec_count_9  <= spec_count_9  + 4'd1;
                        5'd10: spec_count_10 <= spec_count_10 + 4'd1;
                        5'd11: spec_count_11 <= spec_count_11 + 4'd1;
                        5'd12: spec_count_12 <= spec_count_12 + 4'd1;
                        5'd13: spec_count_13 <= spec_count_13 + 4'd1;
                        5'd14: spec_count_14 <= spec_count_14 + 4'd1;
                        5'd15: spec_count_15 <= spec_count_15 + 4'd1;
                        5'd16: spec_count_16 <= spec_count_16 + 4'd1;
                        5'd17: spec_count_17 <= spec_count_17 + 4'd1;
                        5'd18: spec_count_18 <= spec_count_18 + 4'd1;
                        5'd19: spec_count_19 <= spec_count_19 + 4'd1;
                        5'd20: spec_count_20 <= spec_count_20 + 4'd1;
                        5'd21: spec_count_21 <= spec_count_21 + 4'd1;
                        5'd22: spec_count_22 <= spec_count_22 + 4'd1;
                        5'd23: spec_count_23 <= spec_count_23 + 4'd1;
                        5'd24: spec_count_24 <= spec_count_24 + 4'd1;
                        default: ;
                    endcase
                end
                else if (!need_overwrite && !found_empty) begin
                    // ���2�������������need_overwrite=0��û�пղ�λ��
                    // �������䣬�¹�����+1�������ǹ�����-1
                    
                    // �¹�����+1
                    case (spec_idx)
                        5'd0:  spec_count_0  <= spec_count_0  + 4'd1;
                        5'd1:  spec_count_1  <= spec_count_1  + 4'd1;
                        5'd2:  spec_count_2  <= spec_count_2  + 4'd1;
                        5'd3:  spec_count_3  <= spec_count_3  + 4'd1;
                        5'd4:  spec_count_4  <= spec_count_4  + 4'd1;
                        5'd5:  spec_count_5  <= spec_count_5  + 4'd1;
                        5'd6:  spec_count_6  <= spec_count_6  + 4'd1;
                        5'd7:  spec_count_7  <= spec_count_7  + 4'd1;
                        5'd8:  spec_count_8  <= spec_count_8  + 4'd1;
                        5'd9:  spec_count_9  <= spec_count_9  + 4'd1;
                        5'd10: spec_count_10 <= spec_count_10 + 4'd1;
                        5'd11: spec_count_11 <= spec_count_11 + 4'd1;
                        5'd12: spec_count_12 <= spec_count_12 + 4'd1;
                        5'd13: spec_count_13 <= spec_count_13 + 4'd1;
                        5'd14: spec_count_14 <= spec_count_14 + 4'd1;
                        5'd15: spec_count_15 <= spec_count_15 + 4'd1;
                        5'd16: spec_count_16 <= spec_count_16 + 4'd1;
                        5'd17: spec_count_17 <= spec_count_17 + 4'd1;
                        5'd18: spec_count_18 <= spec_count_18 + 4'd1;
                        5'd19: spec_count_19 <= spec_count_19 + 4'd1;
                        5'd20: spec_count_20 <= spec_count_20 + 4'd1;
                        5'd21: spec_count_21 <= spec_count_21 + 4'd1;
                        5'd22: spec_count_22 <= spec_count_22 + 4'd1;
                        5'd23: spec_count_23 <= spec_count_23 + 4'd1;
                        5'd24: spec_count_24 <= spec_count_24 + 4'd1;
                        default: ;
                    endcase
                    
                    // �����ǹ�����-1
                    case (old_spec_idx)
                        5'd0:  spec_count_0  <= spec_count_0  - 4'd1;
                        5'd1:  spec_count_1  <= spec_count_1  - 4'd1;
                        5'd2:  spec_count_2  <= spec_count_2  - 4'd1;
                        5'd3:  spec_count_3  <= spec_count_3  - 4'd1;
                        5'd4:  spec_count_4  <= spec_count_4  - 4'd1;
                        5'd5:  spec_count_5  <= spec_count_5  - 4'd1;
                        5'd6:  spec_count_6  <= spec_count_6  - 4'd1;
                        5'd7:  spec_count_7  <= spec_count_7  - 4'd1;
                        5'd8:  spec_count_8  <= spec_count_8  - 4'd1;
                        5'd9:  spec_count_9  <= spec_count_9  - 4'd1;
                        5'd10: spec_count_10 <= spec_count_10 - 4'd1;
                        5'd11: spec_count_11 <= spec_count_11 - 4'd1;
                        5'd12: spec_count_12 <= spec_count_12 - 4'd1;
                        5'd13: spec_count_13 <= spec_count_13 - 4'd1;
                        5'd14: spec_count_14 <= spec_count_14 - 4'd1;
                        5'd15: spec_count_15 <= spec_count_15 - 4'd1;
                        5'd16: spec_count_16 <= spec_count_16 - 4'd1;
                        5'd17: spec_count_17 <= spec_count_17 - 4'd1;
                        5'd18: spec_count_18 <= spec_count_18 - 4'd1;
                        5'd19: spec_count_19 <= spec_count_19 - 4'd1;
                        5'd20: spec_count_20 <= spec_count_20 - 4'd1;
                        5'd21: spec_count_21 <= spec_count_21 - 4'd1;
                        5'd22: spec_count_22 <= spec_count_22 - 4'd1;
                        5'd23: spec_count_23 <= spec_count_23 - 4'd1;
                        5'd24: spec_count_24 <= spec_count_24 - 4'd1;
                        default: ;
                    endcase
                end
                // ���3������ͬ���need_overwrite=1�������ı��κμ���
            end
            
            //==================================================================
            // ��ȡ������
            //==================================================================
            if (read_en) begin
                read_done <= 1'b1;
                
                case (read_idx)
                    4'd0: begin
                        read_out_m <= mat_m_0; read_out_n <= mat_n_0;
                        read_out_data <= mat_data_0; read_out_id <= mat_id_0;
                        read_valid <= mat_valid_0;
                    end
                    4'd1: begin
                        read_out_m <= mat_m_1; read_out_n <= mat_n_1;
                        read_out_data <= mat_data_1; read_out_id <= mat_id_1;
                        read_valid <= mat_valid_1;
                    end
                    4'd2: begin
                        read_out_m <= mat_m_2; read_out_n <= mat_n_2;
                        read_out_data <= mat_data_2; read_out_id <= mat_id_2;
                        read_valid <= mat_valid_2;
                    end
                    4'd3: begin
                        read_out_m <= mat_m_3; read_out_n <= mat_n_3;
                        read_out_data <= mat_data_3; read_out_id <= mat_id_3;
                        read_valid <= mat_valid_3;
                    end
                    4'd4: begin
                        read_out_m <= mat_m_4; read_out_n <= mat_n_4;
                        read_out_data <= mat_data_4; read_out_id <= mat_id_4;
                        read_valid <= mat_valid_4;
                    end
                    4'd5: begin
                        read_out_m <= mat_m_5; read_out_n <= mat_n_5;
                        read_out_data <= mat_data_5; read_out_id <= mat_id_5;
                        read_valid <= mat_valid_5;
                    end
                    4'd6: begin
                        read_out_m <= mat_m_6; read_out_n <= mat_n_6;
                        read_out_data <= mat_data_6; read_out_id <= mat_id_6;
                        read_valid <= mat_valid_6;
                    end
                    4'd7: begin
                        read_out_m <= mat_m_7; read_out_n <= mat_n_7;
                        read_out_data <= mat_data_7; read_out_id <= mat_id_7;
                        read_valid <= mat_valid_7;
                    end
                    4'd8: begin
                        read_out_m <= mat_m_8; read_out_n <= mat_n_8;
                        read_out_data <= mat_data_8; read_out_id <= mat_id_8;
                        read_valid <= mat_valid_8;
                    end
                    4'd9: begin
                        read_out_m <= mat_m_9; read_out_n <= mat_n_9;
                        read_out_data <= mat_data_9; read_out_id <= mat_id_9;
                        read_valid <= mat_valid_9;
                    end
                    default: begin
                        read_out_m <= 4'd0; read_out_n <= 4'd0;
                        read_out_data <= 200'd0; read_out_id <= 4'd0;
                        read_valid <= 1'b0;
                    end
                endcase
            end
        end
    end

endmodule