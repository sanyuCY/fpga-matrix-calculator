//�����������ģ��
// ģ�鹦�ܣ�����UART��������ľ������ݣ����ά��/Ԫ�غϷ��Լ�⣬����ṹ����������
// ����Vivado 2017����5��5��ά������Ϊ25������4λ�źţ��������˿ڼ�������
module matrix_input(
    input clk,
    input rst_n,// �͵�ƽ��λ��0=��λ��1=����������
    //����UARTģ��
    input [7:0] uart_rx_data, // UART���յĵ��ֽ����ݣ�ASCII�룬8λ��
    input rx_done,      // UART���ֽڽ�����ɱ�־���ߵ�ƽ��Ч������1��ʱ�ӣ�
    // ����FSMģ��
    input [3:0] val_min,
    input [3:0] val_max,
    // ������洢/����ģ��ľ���ά��
    output reg [3:0] mat_m,  // ����������1~5��
    output reg [3:0] mat_n,  // ����������1~5��
    // �����޸ģ�5��5������Ϊ25������4λ�źţ������ά����˿ڣ�
    output reg [3:0] mat_data_00, mat_data_01, mat_data_02, mat_data_03, mat_data_04,
    output reg [3:0] mat_data_10, mat_data_11, mat_data_12, mat_data_13, mat_data_14,
    output reg [3:0] mat_data_20, mat_data_21, mat_data_22, mat_data_23, mat_data_24,
    output reg [3:0] mat_data_30, mat_data_31, mat_data_32, mat_data_33, mat_data_34,
    output reg [3:0] mat_data_40, mat_data_41, mat_data_42, mat_data_43, mat_data_44,
    // �����FSMģ���״̬/�����־
    output reg input_done, // ������ɱ�־���ߵ�ƽ��Ч������1��ʱ�ӣ�
    output reg [2:0] error_type  // �������ͣ�000=�޴�001=ά�ȴ�011=Ԫ��ֵ��
);

// ״̬�����壨��ԭʼ������ȫһ�£�
localparam S_WAIT = 3'b000;     // �ȴ�UART��������
localparam S_PARSE_M = 3'b001;  // ������������m
localparam S_PARSE_N = 3'b010;  // ������������n
localparam S_PARSE_DATA= 3'b011;// ��������Ԫ��
localparam S_CHECK = 3'b100;    // �Ϸ��Լ��
localparam S_DONE = 3'b101;     // ������ɣ�������

// ״̬���Ĵ�������ԭʼ������ȫһ�£�
reg [2:0] curr_state;  // ��ǰ״̬
reg [2:0] next_state;  // ��һ״̬������ʽ״̬����

// ��ʱ�洢�Ĵ������ڲ����ö�ά���飬��Ӱ���߼���д��
reg [3:0] m_temp;      // ������ʱ����
reg [3:0] n_temp;      // ������ʱ����
reg [3:0] data_temp [0:4][0:4]; // Ԫ����ʱ���棨5��5��
reg [4:0] data_cnt;    // Ԫ�ؼ�������0~24��

// ѭ��������������ԭʼ����һ�£�
integer i, j;

// ����1��״̬����ǰ״̬���£�ʱ���ش�����
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        curr_state <= S_WAIT; // ��λ���ʼ״̬���ȴ�
    end else begin
        curr_state <= next_state; // �Ǹ�λʱ����Ϊ��һ״̬
    end
end

// ����2��״̬����һ״̬���㣨����߼���
always @(*) begin
    next_state = curr_state; // Ĭ�ϱ��ֵ�ǰ״̬��������������
    case(curr_state)
        S_WAIT: begin
            // ����������UART�յ���һ���ֽڣ�����m��
            if(rx_done) begin
                next_state = S_PARSE_M;
            end
        end
        S_PARSE_M: begin
            // ����������UART�յ��ڶ����ֽڣ�����n��
            if(rx_done) begin
                next_state = S_PARSE_N;
            end
        end
        S_PARSE_N: begin
            // ����������UART�յ��������ֽڣ���һ��Ԫ�أ�
            if(rx_done) begin
                next_state = S_PARSE_DATA;
            end
        end
        S_PARSE_DATA: begin
            // ����������Ԫ�ؽ�����ɣ��������ﵽm��n-1�����յ����һ��Ԫ��
            if(rx_done && (data_cnt == m_temp * n_temp - 1)) begin
                next_state = S_CHECK;
            end
        end
        S_CHECK: begin
            // �Ϸ��Լ����ɺ󣬽������״̬
            next_state = S_DONE;
        end
        S_DONE: begin
            // ��ɺ�ص��ȴ�״̬��׼����һ�ν���
            next_state = S_WAIT;
        end
        default: begin
            // �쳣״̬�ص��ȴ������³����
            next_state = S_WAIT;
        end
    endcase
end

// ����3��UART�������浽��ʱ�Ĵ�������ԭʼ������ȫһ�£�
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        // ��λ�����������ʱ�Ĵ����ͼ�����
        m_temp <= 4'd0;
        n_temp <= 4'd0;
        data_cnt <= 5'd0;
        // ��ʱ������Ԫ�ظ�λ����ԭʼ����һ�£�
        data_temp[0][0] <= 4'd0;
        data_temp[0][1] <= 4'd0;
        data_temp[0][2] <= 4'd0;
        data_temp[0][3] <= 4'd0;
        data_temp[0][4] <= 4'd0;
        data_temp[1][0] <= 4'd0;
        data_temp[1][1] <= 4'd0;
        data_temp[1][2] <= 4'd0;
        data_temp[1][3] <= 4'd0;
        data_temp[1][4] <= 4'd0;
        data_temp[2][0] <= 4'd0;
        data_temp[2][1] <= 4'd0;
        data_temp[2][2] <= 4'd0;
        data_temp[2][3] <= 4'd0;
        data_temp[2][4] <= 4'd0;
        data_temp[3][0] <= 4'd0;
        data_temp[3][1] <= 4'd0;
        data_temp[3][2] <= 4'd0;
        data_temp[3][3] <= 4'd0;
        data_temp[3][4] <= 4'd0;
        data_temp[4][0] <= 4'd0;
        data_temp[4][1] <= 4'd0;
        data_temp[4][2] <= 4'd0;
        data_temp[4][3] <= 4'd0;
        data_temp[4][4] <= 4'd0;
    end else begin
        case(curr_state)
            S_PARSE_M: begin
                // ASCIIת���֣�ȡ��4λ��0~9��
                if(rx_done) begin
                    m_temp <= uart_rx_data[3:0];
                end
            end
            S_PARSE_N: begin
                // ��������n���������߼�һ��
                if(rx_done) begin
                    n_temp <= uart_rx_data[3:0];
                end
            end
            S_PARSE_DATA: begin
                // ����Ԫ�أ������������洢����ʱ����
                if(rx_done) begin
                    data_temp[data_cnt / n_temp][data_cnt % n_temp] <= uart_rx_data[3:0];
                    data_cnt <= data_cnt + 1'b1; // ����������
                end
            end
            S_DONE: begin
                // ������ɺ����ü�����
                data_cnt <= 5'd0;
            end
            default: begin
                // ����״̬������ʱ�Ĵ�������
                m_temp <= m_temp;
                n_temp <= n_temp;
                data_cnt <= data_cnt;
            end
        endcase
    end
end

// ����4���Ϸ��Լ�� + ��������ֵ�������޸ģ������źŸ�ֵ��
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        // ��λ�������������Ĵ����ͱ�־
        mat_m <= 4'd0;
        mat_n <= 4'd0;
        input_done <= 1'b0;
        error_type <= 3'b000;
        // �����ź���λ��λ����ԭʼ�������鸴λ�߼�һ�£�
        mat_data_00 <= 4'd0; mat_data_01 <= 4'd0; mat_data_02 <= 4'd0; mat_data_03 <= 4'd0; mat_data_04 <= 4'd0;
        mat_data_10 <= 4'd0; mat_data_11 <= 4'd0; mat_data_12 <= 4'd0; mat_data_13 <= 4'd0; mat_data_14 <= 4'd0;
        mat_data_20 <= 4'd0; mat_data_21 <= 4'd0; mat_data_22 <= 4'd0; mat_data_23 <= 4'd0; mat_data_24 <= 4'd0;
        mat_data_30 <= 4'd0; mat_data_31 <= 4'd0; mat_data_32 <= 4'd0; mat_data_33 <= 4'd0; mat_data_34 <= 4'd0;
        mat_data_40 <= 4'd0; mat_data_41 <= 4'd0; mat_data_42 <= 4'd0; mat_data_43 <= 4'd0; mat_data_44 <= 4'd0;
    end else begin
        case(curr_state)
            S_CHECK: begin
                // ��ʼ����������Ϊ�޴�
                error_type <= 3'b000;
                
                // ��һ�������ά�ȺϷ��ԣ�1~5��
                if(m_temp < 4'd1 || m_temp > 4'd5 || n_temp < 4'd1 || n_temp > 4'd5) begin
                    error_type <= 3'b001; // ά�ȴ���
                end else begin
                    // �ڶ��������Ԫ��ֵ�Ϸ��ԣ�val_min~val_max��
                    for(i=0; i<m_temp; i=i+1) begin 
                        for(j=0; j<n_temp; j=j+1) begin 
                            if(data_temp[i][j] < val_min || data_temp[i][j] > val_max) begin
                                error_type <= 3'b011; // Ԫ��ֵ����
                            end
                        end
                    end
                end
            end
            S_DONE: begin
                // ��λ��ɱ�־������FSMģ�������ɣ�
                input_done <= 1'b1;
                
                if(error_type == 3'b000) begin
                    // �޴����������ά�� + �����źŸ�ֵ����ԭʼ����һһ��Ӧ��
                    mat_m <= m_temp;
                    mat_n <= n_temp;
                    // ��Ԫ�ظ�ֵ����ʱ���� �� ��������ź�
                    mat_data_00 <= data_temp[0][0]; mat_data_01 <= data_temp[0][1]; mat_data_02 <= data_temp[0][2]; mat_data_03 <= data_temp[0][3]; mat_data_04 <= data_temp[0][4];
                    mat_data_10 <= data_temp[1][0]; mat_data_11 <= data_temp[1][1]; mat_data_12 <= data_temp[1][2]; mat_data_13 <= data_temp[1][3]; mat_data_14 <= data_temp[1][4];
                    mat_data_20 <= data_temp[2][0]; mat_data_21 <= data_temp[2][1]; mat_data_22 <= data_temp[2][2]; mat_data_23 <= data_temp[2][3]; mat_data_24 <= data_temp[2][4];
                    mat_data_30 <= data_temp[3][0]; mat_data_31 <= data_temp[3][1]; mat_data_32 <= data_temp[3][2]; mat_data_33 <= data_temp[3][3]; mat_data_34 <= data_temp[3][4];
                    mat_data_40 <= data_temp[4][0]; mat_data_41 <= data_temp[4][1]; mat_data_42 <= data_temp[4][2]; mat_data_43 <= data_temp[4][3]; mat_data_44 <= data_temp[4][4];
                end else begin
                    // �д������������������������Ч���ݣ�
                    mat_m <= 4'd0;
                    mat_n <= 4'd0;
                    mat_data_00 <= 4'd0; mat_data_01 <= 4'd0; mat_data_02 <= 4'd0; mat_data_03 <= 4'd0; mat_data_04 <= 4'd0;
                    mat_data_10 <= 4'd0; mat_data_11 <= 4'd0; mat_data_12 <= 4'd0; mat_data_13 <= 4'd0; mat_data_14 <= 4'd0;
                    mat_data_20 <= 4'd0; mat_data_21 <= 4'd0; mat_data_22 <= 4'd0; mat_data_23 <= 4'd0; mat_data_24 <= 4'd0;
                    mat_data_30 <= 4'd0; mat_data_31 <= 4'd0; mat_data_32 <= 4'd0; mat_data_33 <= 4'd0; mat_data_34 <= 4'd0;
                    mat_data_40 <= 4'd0; mat_data_41 <= 4'd0; mat_data_42 <= 4'd0; mat_data_43 <= 4'd0; mat_data_44 <= 4'd0;
                end
            end
            default: begin
                // ����״̬�������ɱ�־�����ִ�������
                input_done <= 1'b0;
                error_type <= error_type;
            end
        endcase
    end
end

endmodule