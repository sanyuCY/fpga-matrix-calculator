module matrix_input(
    input clk,
    input rst_n,
    input [7:0] uart_rx_data,
    input rx_done,
    input [3:0] val_min,
    input [3:0] val_max,
    output reg [3:0] mat_m,
    output reg [3:0] mat_n,
    output reg [3:0] mat_data_00, mat_data_01,
    output reg input_done,
    output reg [2:0] error_type
);

// �����������źţ�ȥ���޹ص�mat_data_xx�����ٸ���
reg [1:0] step;       // ���ղ��裺0=����m��1=����n��2=����Ԫ�أ�3=���
reg [3:0] m_cache;    // ����m
reg [3:0] n_cache;    // ����n
reg [3:0] elem1;      // �����һ��Ԫ�أ�0,0��
reg [3:0] elem2;      // ����ڶ���Ԫ�أ�0,1��
reg [1:0] elem_cnt;   // Ԫ�ؼ���

// ����1���ֽ׶ν���m/n/Ԫ�أ��޳��㣬�޼���������
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        step <= 2'd0;
        m_cache <= 4'd0;
        n_cache <= 4'd0;
        elem1 <= 4'd0;
        elem2 <= 4'd0;
        elem_cnt <= 2'd0;
    end else begin
        if(rx_done) begin
            case(step)
                2'd0: begin // ����m
                    m_cache <= uart_rx_data[3:0];
                    step <= 2'd1;
                end
                2'd1: begin // ����n
                    n_cache <= uart_rx_data[3:0];
                    step <= 2'd2;
                end
                2'd2: begin // ����Ԫ�أ���2x2��
                    if(elem_cnt == 2'd0) begin
                        elem1 <= uart_rx_data[3:0]; // ��һ��Ԫ��
                        elem_cnt <= 2'd1;
                    end else if(elem_cnt == 2'd1) begin
                        elem2 <= uart_rx_data[3:0]; // �ڶ���Ԫ��
                        step <= 2'd3; // �������
                    end
                end
            endcase
        end
    end
end

// ����2��ֱ�Ӹ�ֵ������޸���������ǿ����Ч��
always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        mat_m <= 4'd0;
        mat_n <= 4'd0;
        mat_data_00 <= 4'd0;
        mat_data_01 <= 4'd0;
        input_done <= 1'b0;
        error_type <= 3'b000;
    end else begin
        // Ĭ��ֵ
        input_done <= 1'b0;
        error_type <= 3'b000;

        // ����3=��ɣ���ʼ��ֵ
        if(step == 2'd3) begin
            input_done <= 1'b1;
            // ά�ȼ��
            if(m_cache < 1 || m_cache > 5 || n_cache < 1 || n_cache > 5) begin
                error_type <= 3'b001;
                mat_m <= 4'd0;
                mat_n <= 4'd0;
                mat_data_00 <= 4'd0;
                mat_data_01 <= 4'd0;
            end else begin
                // Ԫ�ؼ��
                if(elem1 < val_min || elem1 > val_max || elem2 < val_min || elem2 > val_max) begin
                    error_type <= 3'b011;
                    mat_m <= 4'd0;
                    mat_n <= 4'd0;
                    mat_data_00 <= 4'd0;
                    mat_data_01 <= 4'd0;
                end else begin
                    // ǿ�Ƹ�ֵ��100%��Ч
                    mat_m <= m_cache;
                    mat_n <= n_cache;
                    mat_data_00 <= elem1;
                    mat_data_01 <= elem2;
                end
            end
        end
    end
end

endmodule